// write your module here
module isodd (
    input [3:0] a,
    output x
);
assign x = a[0];
endmodule